// Benchmark "rand11" written by ABC on Mon Mar  7 02:11:18 2016

module ckt_org ( 
    i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i10,
    f  );
  input  i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i10;
  output f;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
    n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713;
  assign n13 = ~i09 & i10;
  assign n14 = i09 & ~i10;
  assign n15 = ~n13 & ~n14;
  assign n16 = i03 & i06;
  assign n17 = ~i07 & i08;
  assign n18 = n16 & n17;
  assign n19 = ~i03 & ~i06;
  assign n20 = i07 & ~i08;
  assign n21 = n19 & n20;
  assign n22 = ~n18 & ~n21;
  assign n23 = i00 & ~n22;
  assign n24 = ~i06 & i07;
  assign n25 = i03 & n24;
  assign n26 = i06 & ~i07;
  assign n27 = ~i03 & n26;
  assign n28 = ~n25 & ~n27;
  assign n29 = ~i08 & ~n28;
  assign n30 = ~i00 & n29;
  assign n31 = ~n23 & ~n30;
  assign n32 = ~i02 & ~n31;
  assign n33 = ~i07 & ~i08;
  assign n34 = ~i03 & n33;
  assign n35 = i02 & n34;
  assign n36 = ~i00 & n35;
  assign n37 = ~n32 & ~n36;
  assign n38 = i01 & i04;
  assign n39 = ~i01 & ~i04;
  assign n40 = ~n38 & ~n39;
  assign n41 = ~n37 & ~n40;
  assign n42 = ~i01 & i04;
  assign n43 = i01 & ~i04;
  assign n44 = ~n42 & ~n43;
  assign n45 = ~i06 & ~i08;
  assign n46 = ~i00 & n45;
  assign n47 = i00 & ~i03;
  assign n48 = i06 & i08;
  assign n49 = n47 & n48;
  assign n50 = ~n46 & ~n49;
  assign n51 = i07 & ~n50;
  assign n52 = i03 & n33;
  assign n53 = ~i00 & n52;
  assign n54 = ~n51 & ~n53;
  assign n55 = ~n44 & ~n54;
  assign n56 = ~i04 & i08;
  assign n57 = i03 & n56;
  assign n58 = i04 & ~i08;
  assign n59 = ~i03 & n58;
  assign n60 = ~n57 & ~n59;
  assign n61 = ~i01 & ~n60;
  assign n62 = i03 & ~i04;
  assign n63 = i03 & ~n62;
  assign n64 = i08 & ~n63;
  assign n65 = i01 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~i00 & ~n66;
  assign n68 = ~i03 & ~i08;
  assign n69 = ~i03 & ~n68;
  assign n70 = ~i04 & ~n69;
  assign n71 = i01 & n70;
  assign n72 = i00 & n71;
  assign n73 = ~n67 & ~n72;
  assign n74 = ~i07 & ~n73;
  assign n75 = ~i00 & i03;
  assign n76 = ~i00 & ~n75;
  assign n77 = i08 & ~n76;
  assign n78 = i07 & n77;
  assign n79 = i04 & n78;
  assign n80 = i01 & n79;
  assign n81 = ~n74 & ~n80;
  assign n82 = ~i06 & ~n81;
  assign n83 = ~i03 & i08;
  assign n84 = i03 & ~i08;
  assign n85 = ~n83 & ~n84;
  assign n86 = ~i07 & ~n85;
  assign n87 = i06 & n86;
  assign n88 = i04 & n87;
  assign n89 = i01 & n88;
  assign n90 = ~i00 & n89;
  assign n91 = ~n82 & ~n90;
  assign n92 = ~n55 & n91;
  assign n93 = i02 & ~n92;
  assign n94 = i00 & n24;
  assign n95 = ~i00 & n26;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~i01 & ~i03;
  assign n98 = i04 & i08;
  assign n99 = n97 & n98;
  assign n100 = i01 & i03;
  assign n101 = ~i04 & ~i08;
  assign n102 = n100 & n101;
  assign n103 = ~n99 & ~n102;
  assign n104 = ~n96 & ~n103;
  assign n105 = ~i00 & ~i07;
  assign n106 = ~i00 & ~n105;
  assign n107 = ~i03 & ~i04;
  assign n108 = ~i06 & i08;
  assign n109 = n107 & n108;
  assign n110 = i03 & i04;
  assign n111 = i06 & ~i08;
  assign n112 = n110 & n111;
  assign n113 = ~n109 & ~n112;
  assign n114 = ~n106 & ~n113;
  assign n115 = i03 & i07;
  assign n116 = ~i03 & ~i07;
  assign n117 = ~n115 & ~n116;
  assign n118 = i00 & ~n117;
  assign n119 = ~i03 & i07;
  assign n120 = ~i00 & n119;
  assign n121 = ~n118 & ~n120;
  assign n122 = i08 & ~n121;
  assign n123 = ~i00 & ~i03;
  assign n124 = n20 & n123;
  assign n125 = ~n122 & ~n124;
  assign n126 = i06 & ~n125;
  assign n127 = i03 & ~i07;
  assign n128 = ~i03 & n20;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~i06 & ~n129;
  assign n131 = ~i00 & n130;
  assign n132 = ~n126 & ~n131;
  assign n133 = i04 & ~n132;
  assign n134 = ~i00 & n107;
  assign n135 = ~i06 & n33;
  assign n136 = n134 & n135;
  assign n137 = ~n133 & ~n136;
  assign n138 = ~n114 & n137;
  assign n139 = i01 & ~n138;
  assign n140 = ~n108 & ~n111;
  assign n141 = ~i00 & ~n140;
  assign n142 = i00 & n48;
  assign n143 = ~n141 & ~n142;
  assign n144 = i07 & ~n143;
  assign n145 = i00 & n33;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~i03 & ~n146;
  assign n148 = i06 & i07;
  assign n149 = ~i06 & ~i07;
  assign n150 = ~n148 & ~n149;
  assign n151 = i00 & ~n150;
  assign n152 = ~i00 & n148;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~i08 & ~n153;
  assign n155 = i03 & n154;
  assign n156 = ~n147 & ~n155;
  assign n157 = i04 & ~n156;
  assign n158 = ~i01 & n157;
  assign n159 = ~n139 & ~n158;
  assign n160 = ~n104 & n159;
  assign n161 = ~i02 & ~n160;
  assign n162 = ~n93 & ~n161;
  assign n163 = ~n41 & n162;
  assign n164 = ~i05 & ~n163;
  assign n165 = i03 & n148;
  assign n166 = ~i03 & n149;
  assign n167 = ~n165 & ~n166;
  assign n168 = i02 & ~n167;
  assign n169 = i06 & ~n26;
  assign n170 = ~i03 & ~n169;
  assign n171 = i03 & n149;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~i02 & ~n172;
  assign n174 = ~n168 & ~n173;
  assign n175 = ~i04 & ~n174;
  assign n176 = i02 & ~i07;
  assign n177 = i02 & ~n176;
  assign n178 = i06 & ~n177;
  assign n179 = i04 & n178;
  assign n180 = ~i03 & n179;
  assign n181 = ~n175 & ~n180;
  assign n182 = ~i08 & ~n181;
  assign n183 = ~i03 & ~n119;
  assign n184 = ~i06 & ~n183;
  assign n185 = ~i03 & n148;
  assign n186 = ~n184 & ~n185;
  assign n187 = i04 & ~n186;
  assign n188 = ~i04 & ~n150;
  assign n189 = ~i03 & n188;
  assign n190 = ~n187 & ~n189;
  assign n191 = i02 & ~n190;
  assign n192 = ~n27 & ~n115;
  assign n193 = i04 & ~n192;
  assign n194 = ~i02 & n193;
  assign n195 = ~n191 & ~n194;
  assign n196 = i08 & ~n195;
  assign n197 = ~n182 & ~n196;
  assign n198 = ~i00 & ~n197;
  assign n199 = i02 & i07;
  assign n200 = ~i02 & ~i07;
  assign n201 = ~n199 & ~n200;
  assign n202 = ~i03 & i06;
  assign n203 = i04 & ~i06;
  assign n204 = i03 & n203;
  assign n205 = ~n202 & ~n204;
  assign n206 = ~n201 & ~n205;
  assign n207 = ~n16 & ~n19;
  assign n208 = i02 & ~n207;
  assign n209 = ~i02 & n16;
  assign n210 = ~n208 & ~n209;
  assign n211 = ~i07 & ~n210;
  assign n212 = i04 & n211;
  assign n213 = ~n206 & ~n212;
  assign n214 = ~i08 & ~n213;
  assign n215 = ~i02 & n24;
  assign n216 = i02 & n26;
  assign n217 = ~n215 & ~n216;
  assign n218 = i02 & ~i04;
  assign n219 = n24 & n218;
  assign n220 = n217 & ~n219;
  assign n221 = i03 & ~n220;
  assign n222 = i04 & n149;
  assign n223 = ~n188 & ~n222;
  assign n224 = ~i03 & ~n223;
  assign n225 = ~i02 & n224;
  assign n226 = ~n221 & ~n225;
  assign n227 = i08 & ~n226;
  assign n228 = ~n214 & ~n227;
  assign n229 = i00 & ~n228;
  assign n230 = ~n198 & ~n229;
  assign n231 = i01 & ~n230;
  assign n232 = i07 & i08;
  assign n233 = i06 & n232;
  assign n234 = ~n135 & ~n233;
  assign n235 = ~i03 & i04;
  assign n236 = ~n62 & ~n235;
  assign n237 = ~i00 & ~n236;
  assign n238 = i00 & n62;
  assign n239 = ~n237 & ~n238;
  assign n240 = ~n234 & ~n239;
  assign n241 = ~i04 & n108;
  assign n242 = i04 & n111;
  assign n243 = ~n241 & ~n242;
  assign n244 = i03 & ~n243;
  assign n245 = ~i04 & n48;
  assign n246 = ~n58 & ~n245;
  assign n247 = ~i03 & ~n246;
  assign n248 = ~n244 & ~n247;
  assign n249 = i07 & ~n248;
  assign n250 = n135 & n235;
  assign n251 = ~n249 & ~n250;
  assign n252 = i00 & ~n251;
  assign n253 = ~i04 & ~n56;
  assign n254 = ~i07 & ~n253;
  assign n255 = ~i04 & n232;
  assign n256 = ~n254 & ~n255;
  assign n257 = i06 & ~n256;
  assign n258 = ~i03 & n257;
  assign n259 = ~i00 & n258;
  assign n260 = ~n252 & ~n259;
  assign n261 = ~n240 & n260;
  assign n262 = ~i02 & ~n261;
  assign n263 = i04 & n232;
  assign n264 = ~i04 & n33;
  assign n265 = ~n263 & ~n264;
  assign n266 = i03 & ~n265;
  assign n267 = n20 & n107;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~i06 & ~n268;
  assign n270 = n107 & n233;
  assign n271 = ~n269 & ~n270;
  assign n272 = i04 & i06;
  assign n273 = ~i04 & ~i06;
  assign n274 = ~n272 & ~n273;
  assign n275 = i03 & ~n274;
  assign n276 = ~i03 & n272;
  assign n277 = ~n275 & ~n276;
  assign n278 = ~i00 & n17;
  assign n279 = i00 & n20;
  assign n280 = ~n278 & ~n279;
  assign n281 = ~n277 & ~n280;
  assign n282 = i04 & ~n234;
  assign n283 = i03 & n282;
  assign n284 = n107 & n135;
  assign n285 = ~n283 & ~n284;
  assign n286 = i00 & ~n285;
  assign n287 = ~n281 & ~n286;
  assign n288 = n271 & n287;
  assign n289 = i02 & ~n288;
  assign n290 = ~n262 & ~n289;
  assign n291 = ~i01 & ~n290;
  assign n292 = ~n231 & ~n291;
  assign n293 = i05 & ~n292;
  assign n294 = ~n164 & ~n293;
  assign n295 = ~n15 & ~n294;
  assign n296 = i04 & n45;
  assign n297 = ~n245 & ~n296;
  assign n298 = i09 & i10;
  assign n299 = i02 & n298;
  assign n300 = ~i09 & ~i10;
  assign n301 = ~i02 & n300;
  assign n302 = ~n299 & ~n301;
  assign n303 = ~i05 & ~n302;
  assign n304 = i00 & n303;
  assign n305 = ~i00 & ~i02;
  assign n306 = i05 & n14;
  assign n307 = n305 & n306;
  assign n308 = ~n304 & ~n307;
  assign n309 = i01 & ~n308;
  assign n310 = ~i01 & i02;
  assign n311 = ~i00 & n310;
  assign n312 = i05 & n300;
  assign n313 = n311 & n312;
  assign n314 = ~n309 & ~n313;
  assign n315 = n200 & n298;
  assign n316 = n199 & n300;
  assign n317 = ~n315 & ~n316;
  assign n318 = i05 & ~n317;
  assign n319 = i00 & n318;
  assign n320 = ~i02 & i07;
  assign n321 = n298 & n320;
  assign n322 = n176 & n300;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~i05 & ~n323;
  assign n325 = ~i00 & n324;
  assign n326 = ~n319 & ~n325;
  assign n327 = i05 & i09;
  assign n328 = ~i05 & ~i09;
  assign n329 = ~n327 & ~n328;
  assign n330 = i10 & ~n329;
  assign n331 = i02 & n330;
  assign n332 = i00 & n331;
  assign n333 = n305 & n312;
  assign n334 = ~n332 & ~n333;
  assign n335 = i07 & ~n334;
  assign n336 = ~i07 & ~i09;
  assign n337 = ~i05 & n336;
  assign n338 = ~i02 & n337;
  assign n339 = ~i00 & n338;
  assign n340 = ~n335 & ~n339;
  assign n341 = ~i01 & ~n340;
  assign n342 = i07 & i10;
  assign n343 = ~i07 & ~i10;
  assign n344 = ~n342 & ~n343;
  assign n345 = ~i09 & ~n344;
  assign n346 = i05 & n345;
  assign n347 = i02 & n346;
  assign n348 = i01 & n347;
  assign n349 = ~i00 & n348;
  assign n350 = ~n341 & ~n349;
  assign n351 = n326 & n350;
  assign n352 = n314 & n351;
  assign n353 = i03 & ~n352;
  assign n354 = i05 & i07;
  assign n355 = ~i05 & ~i07;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n298 & ~n300;
  assign n358 = i00 & ~n357;
  assign n359 = ~i00 & n298;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~i01 & ~n360;
  assign n362 = ~i00 & i01;
  assign n363 = n300 & n362;
  assign n364 = ~n361 & ~n363;
  assign n365 = ~n356 & ~n364;
  assign n366 = ~i01 & ~i05;
  assign n367 = ~i00 & n366;
  assign n368 = i07 & n298;
  assign n369 = n367 & n368;
  assign n370 = ~n365 & ~n369;
  assign n371 = i02 & ~n370;
  assign n372 = i01 & i05;
  assign n373 = n298 & n372;
  assign n374 = n300 & n366;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~i07 & n13;
  assign n377 = i07 & n14;
  assign n378 = ~n376 & ~n377;
  assign n379 = i05 & ~n378;
  assign n380 = ~i05 & i07;
  assign n381 = n298 & n380;
  assign n382 = ~n379 & ~n381;
  assign n383 = i01 & ~n382;
  assign n384 = n375 & ~n383;
  assign n385 = ~i00 & ~n384;
  assign n386 = i01 & ~i05;
  assign n387 = i00 & n386;
  assign n388 = ~i07 & n298;
  assign n389 = n387 & n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = ~i02 & ~n390;
  assign n392 = ~n371 & ~n391;
  assign n393 = ~i03 & ~n392;
  assign n394 = ~n353 & ~n393;
  assign n395 = ~n297 & ~n394;
  assign n396 = ~i04 & i07;
  assign n397 = ~i08 & n298;
  assign n398 = n396 & n397;
  assign n399 = i04 & ~i07;
  assign n400 = i08 & n300;
  assign n401 = n399 & n400;
  assign n402 = ~n398 & ~n401;
  assign n403 = ~i02 & i06;
  assign n404 = ~i00 & n403;
  assign n405 = i02 & ~i06;
  assign n406 = i00 & n405;
  assign n407 = ~n404 & ~n406;
  assign n408 = ~n402 & ~n407;
  assign n409 = i00 & ~i08;
  assign n410 = ~i00 & n108;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~i09 & ~n411;
  assign n413 = ~i04 & n412;
  assign n414 = ~i00 & i04;
  assign n415 = i08 & i09;
  assign n416 = i06 & n415;
  assign n417 = n414 & n416;
  assign n418 = ~n413 & ~n417;
  assign n419 = ~i10 & ~n418;
  assign n420 = ~i07 & n419;
  assign n421 = ~i00 & n272;
  assign n422 = n20 & n298;
  assign n423 = n421 & n422;
  assign n424 = ~n420 & ~n423;
  assign n425 = ~i02 & ~n424;
  assign n426 = ~n408 & ~n425;
  assign n427 = i03 & ~n426;
  assign n428 = ~i04 & n298;
  assign n429 = i04 & n300;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~i02 & ~n430;
  assign n432 = i00 & n431;
  assign n433 = ~i00 & i02;
  assign n434 = i04 & n298;
  assign n435 = n433 & n434;
  assign n436 = ~n432 & ~n435;
  assign n437 = ~i07 & ~n436;
  assign n438 = i07 & ~n357;
  assign n439 = ~i04 & n438;
  assign n440 = i02 & n439;
  assign n441 = ~i00 & n440;
  assign n442 = ~n437 & ~n441;
  assign n443 = ~i06 & ~n442;
  assign n444 = ~i02 & i04;
  assign n445 = ~i00 & n444;
  assign n446 = n148 & n298;
  assign n447 = n445 & n446;
  assign n448 = ~n443 & ~n447;
  assign n449 = i08 & ~n448;
  assign n450 = n272 & n305;
  assign n451 = n20 & n300;
  assign n452 = n450 & n451;
  assign n453 = ~n449 & ~n452;
  assign n454 = ~i03 & ~n453;
  assign n455 = ~n427 & ~n454;
  assign n456 = ~n17 & ~n20;
  assign n457 = ~n403 & ~n405;
  assign n458 = i10 & ~n457;
  assign n459 = i01 & n458;
  assign n460 = ~i06 & ~i10;
  assign n461 = n310 & n460;
  assign n462 = ~n459 & ~n461;
  assign n463 = ~i03 & ~n462;
  assign n464 = i01 & ~i02;
  assign n465 = i06 & i10;
  assign n466 = i03 & n465;
  assign n467 = n464 & n466;
  assign n468 = ~n463 & ~n467;
  assign n469 = i04 & ~n468;
  assign n470 = i00 & n469;
  assign n471 = i01 & i02;
  assign n472 = ~i00 & n471;
  assign n473 = i06 & ~i10;
  assign n474 = n107 & n473;
  assign n475 = n472 & n474;
  assign n476 = ~n470 & ~n475;
  assign n477 = ~n456 & ~n476;
  assign n478 = ~n97 & ~n100;
  assign n479 = i08 & i10;
  assign n480 = n399 & n479;
  assign n481 = ~i08 & ~i10;
  assign n482 = n396 & n481;
  assign n483 = ~n480 & ~n482;
  assign n484 = i06 & ~n483;
  assign n485 = i02 & n484;
  assign n486 = ~i02 & n273;
  assign n487 = ~i08 & i10;
  assign n488 = ~i07 & n487;
  assign n489 = n486 & n488;
  assign n490 = ~n485 & ~n489;
  assign n491 = i00 & ~n490;
  assign n492 = ~i00 & n218;
  assign n493 = i08 & ~i10;
  assign n494 = n24 & n493;
  assign n495 = n492 & n494;
  assign n496 = ~n491 & ~n495;
  assign n497 = ~n478 & ~n496;
  assign n498 = ~i03 & n396;
  assign n499 = i03 & n399;
  assign n500 = ~n498 & ~n499;
  assign n501 = i02 & n108;
  assign n502 = n403 & n487;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n500 & ~n503;
  assign n505 = i04 & n24;
  assign n506 = ~i04 & n26;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~i03 & ~n507;
  assign n509 = i02 & n508;
  assign n510 = ~i02 & i03;
  assign n511 = n505 & n510;
  assign n512 = ~n509 & ~n511;
  assign n513 = i10 & ~n512;
  assign n514 = ~i02 & n62;
  assign n515 = i06 & n343;
  assign n516 = n514 & n515;
  assign n517 = ~n513 & ~n516;
  assign n518 = i08 & ~n517;
  assign n519 = i02 & n107;
  assign n520 = n24 & n487;
  assign n521 = n519 & n520;
  assign n522 = ~n518 & ~n521;
  assign n523 = ~n504 & n522;
  assign n524 = i01 & ~n523;
  assign n525 = i04 & n108;
  assign n526 = ~i04 & n111;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~i02 & ~n527;
  assign n529 = n108 & n218;
  assign n530 = ~n528 & ~n529;
  assign n531 = i03 & ~n530;
  assign n532 = ~i03 & n111;
  assign n533 = i02 & n532;
  assign n534 = ~n531 & ~n533;
  assign n535 = ~i07 & ~n534;
  assign n536 = i02 & n98;
  assign n537 = ~i02 & n101;
  assign n538 = ~n536 & ~n537;
  assign n539 = i07 & ~n538;
  assign n540 = ~i06 & n539;
  assign n541 = i03 & n540;
  assign n542 = ~n535 & ~n541;
  assign n543 = i10 & ~n542;
  assign n544 = ~i01 & n543;
  assign n545 = ~n524 & ~n544;
  assign n546 = i00 & ~n545;
  assign n547 = i03 & i08;
  assign n548 = ~n68 & ~n547;
  assign n549 = ~i07 & ~n548;
  assign n550 = i02 & n549;
  assign n551 = ~i02 & ~i03;
  assign n552 = n232 & n551;
  assign n553 = ~n550 & ~n552;
  assign n554 = i01 & ~n553;
  assign n555 = ~i02 & ~n320;
  assign n556 = i03 & ~n555;
  assign n557 = ~i02 & n116;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~i08 & ~n558;
  assign n560 = ~i01 & n559;
  assign n561 = ~n554 & ~n560;
  assign n562 = ~i06 & ~n561;
  assign n563 = ~i02 & n86;
  assign n564 = i02 & i03;
  assign n565 = n20 & n564;
  assign n566 = ~n563 & ~n565;
  assign n567 = i06 & ~n566;
  assign n568 = ~i01 & n567;
  assign n569 = ~n562 & ~n568;
  assign n570 = ~i04 & ~n569;
  assign n571 = i01 & ~n150;
  assign n572 = ~i01 & n24;
  assign n573 = ~n571 & ~n572;
  assign n574 = i03 & ~n573;
  assign n575 = n26 & n97;
  assign n576 = ~n574 & ~n575;
  assign n577 = i08 & ~n576;
  assign n578 = i06 & n33;
  assign n579 = n97 & n578;
  assign n580 = ~n577 & ~n579;
  assign n581 = i04 & ~n580;
  assign n582 = i02 & n581;
  assign n583 = ~n570 & ~n582;
  assign n584 = i10 & ~n583;
  assign n585 = ~i00 & n584;
  assign n586 = ~n546 & ~n585;
  assign n587 = ~n497 & n586;
  assign n588 = ~n477 & n587;
  assign n589 = i09 & ~n588;
  assign n590 = ~i06 & i10;
  assign n591 = i03 & n590;
  assign n592 = ~i03 & n473;
  assign n593 = ~n591 & ~n592;
  assign n594 = i00 & ~n593;
  assign n595 = ~i10 & ~n207;
  assign n596 = ~i00 & n595;
  assign n597 = ~n594 & ~n596;
  assign n598 = i04 & ~n597;
  assign n599 = ~i00 & n590;
  assign n600 = i00 & n473;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~i04 & ~n601;
  assign n603 = i03 & n602;
  assign n604 = ~n598 & ~n603;
  assign n605 = i07 & ~n604;
  assign n606 = i00 & ~i04;
  assign n607 = ~i00 & n203;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~i10 & ~n608;
  assign n610 = ~i07 & n609;
  assign n611 = ~i03 & n610;
  assign n612 = ~n605 & ~n611;
  assign n613 = i01 & ~n612;
  assign n614 = ~i10 & ~n500;
  assign n615 = i00 & n614;
  assign n616 = ~i07 & i10;
  assign n617 = ~i04 & n616;
  assign n618 = n123 & n617;
  assign n619 = ~n615 & ~n618;
  assign n620 = ~i06 & ~n619;
  assign n621 = ~i07 & ~n616;
  assign n622 = i06 & ~n621;
  assign n623 = ~i04 & n622;
  assign n624 = i03 & n623;
  assign n625 = ~i00 & n624;
  assign n626 = ~n620 & ~n625;
  assign n627 = ~i01 & ~n626;
  assign n628 = ~n613 & ~n627;
  assign n629 = ~i08 & ~n628;
  assign n630 = n75 & n465;
  assign n631 = ~n594 & ~n630;
  assign n632 = ~i01 & ~n631;
  assign n633 = n362 & n592;
  assign n634 = ~n632 & ~n633;
  assign n635 = i04 & ~n634;
  assign n636 = ~i01 & i10;
  assign n637 = i01 & ~i10;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~i06 & ~n638;
  assign n640 = ~i04 & n639;
  assign n641 = ~i03 & n640;
  assign n642 = i00 & n641;
  assign n643 = ~n635 & ~n642;
  assign n644 = i07 & ~n643;
  assign n645 = ~i04 & i06;
  assign n646 = i01 & n645;
  assign n647 = ~i01 & n203;
  assign n648 = ~n646 & ~n647;
  assign n649 = i10 & ~n648;
  assign n650 = ~i07 & n649;
  assign n651 = ~i03 & n650;
  assign n652 = i00 & n651;
  assign n653 = ~n644 & ~n652;
  assign n654 = i08 & ~n653;
  assign n655 = ~n629 & ~n654;
  assign n656 = ~i02 & ~n655;
  assign n657 = i00 & ~n207;
  assign n658 = ~n75 & ~n657;
  assign n659 = ~i01 & ~n658;
  assign n660 = n202 & n362;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~i10 & ~n661;
  assign n663 = n362 & n466;
  assign n664 = ~n662 & ~n663;
  assign n665 = i08 & ~n664;
  assign n666 = ~i03 & i10;
  assign n667 = ~i01 & n666;
  assign n668 = i03 & ~i10;
  assign n669 = i01 & n668;
  assign n670 = ~n667 & ~n669;
  assign n671 = ~i08 & ~n670;
  assign n672 = i06 & n671;
  assign n673 = i00 & n672;
  assign n674 = ~n665 & ~n673;
  assign n675 = ~i07 & ~n674;
  assign n676 = i00 & n493;
  assign n677 = n123 & n487;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~i06 & ~n678;
  assign n680 = i01 & n679;
  assign n681 = ~i01 & i03;
  assign n682 = ~i00 & n681;
  assign n683 = i06 & n479;
  assign n684 = n682 & n683;
  assign n685 = ~n680 & ~n684;
  assign n686 = i07 & ~n685;
  assign n687 = ~n675 & ~n686;
  assign n688 = i04 & ~n687;
  assign n689 = i01 & i06;
  assign n690 = ~i01 & ~i06;
  assign n691 = ~n689 & ~n690;
  assign n692 = i08 & ~n691;
  assign n693 = i07 & n692;
  assign n694 = i00 & n693;
  assign n695 = n135 & n362;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~i03 & ~n696;
  assign n698 = ~i01 & i07;
  assign n699 = i01 & ~i07;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~i08 & ~n700;
  assign n702 = i06 & n701;
  assign n703 = i03 & n702;
  assign n704 = ~i00 & n703;
  assign n705 = ~n697 & ~n704;
  assign n706 = ~i10 & ~n705;
  assign n707 = n17 & n689;
  assign n708 = n20 & n690;
  assign n709 = ~n707 & ~n708;
  assign n710 = i10 & ~n709;
  assign n711 = i03 & n710;
  assign n712 = ~i00 & n711;
  assign n713 = ~n706 & ~n712;
  assign n714 = ~i04 & ~n713;
  assign n715 = ~n688 & ~n714;
  assign n716 = i02 & ~n715;
  assign n717 = ~n656 & ~n716;
  assign n718 = ~i09 & ~n717;
  assign n719 = ~n589 & ~n718;
  assign n720 = n455 & n719;
  assign n721 = ~i02 & i08;
  assign n722 = i02 & ~i08;
  assign n723 = ~n721 & ~n722;
  assign n724 = i00 & n26;
  assign n725 = ~i00 & ~i06;
  assign n726 = i07 & ~i09;
  assign n727 = n725 & n726;
  assign n728 = ~n724 & ~n727;
  assign n729 = i03 & ~n728;
  assign n730 = ~i07 & i09;
  assign n731 = ~i06 & n730;
  assign n732 = n123 & n731;
  assign n733 = ~n729 & ~n732;
  assign n734 = i05 & ~n733;
  assign n735 = i03 & ~i05;
  assign n736 = i00 & n735;
  assign n737 = i07 & i09;
  assign n738 = i06 & n737;
  assign n739 = n736 & n738;
  assign n740 = ~n734 & ~n739;
  assign n741 = i10 & ~n740;
  assign n742 = ~i06 & n300;
  assign n743 = ~i05 & n742;
  assign n744 = i03 & n743;
  assign n745 = i00 & n744;
  assign n746 = ~n741 & ~n745;
  assign n747 = i04 & ~n746;
  assign n748 = i10 & ~n207;
  assign n749 = i00 & n748;
  assign n750 = n123 & n473;
  assign n751 = ~n749 & ~n750;
  assign n752 = i07 & ~n751;
  assign n753 = ~i05 & n752;
  assign n754 = ~i03 & i05;
  assign n755 = ~i00 & n754;
  assign n756 = ~i06 & n343;
  assign n757 = n755 & n756;
  assign n758 = ~n753 & ~n757;
  assign n759 = i09 & ~n758;
  assign n760 = i07 & n300;
  assign n761 = i05 & n760;
  assign n762 = i03 & n761;
  assign n763 = i00 & n762;
  assign n764 = ~n759 & ~n763;
  assign n765 = ~i04 & ~n764;
  assign n766 = ~n747 & ~n765;
  assign n767 = ~i01 & ~n766;
  assign n768 = i05 & i10;
  assign n769 = ~i05 & ~i10;
  assign n770 = ~n768 & ~n769;
  assign n771 = ~i09 & ~n770;
  assign n772 = ~i06 & n771;
  assign n773 = i00 & n772;
  assign n774 = ~i00 & ~i05;
  assign n775 = i06 & n298;
  assign n776 = n774 & n775;
  assign n777 = ~n773 & ~n776;
  assign n778 = ~i07 & ~n777;
  assign n779 = i06 & n438;
  assign n780 = ~i05 & n779;
  assign n781 = ~i00 & n780;
  assign n782 = ~n778 & ~n781;
  assign n783 = i04 & ~n782;
  assign n784 = ~i05 & i06;
  assign n785 = i07 & n13;
  assign n786 = n784 & n785;
  assign n787 = i05 & ~i06;
  assign n788 = ~i07 & n14;
  assign n789 = n787 & n788;
  assign n790 = ~n786 & ~n789;
  assign n791 = ~i00 & ~n790;
  assign n792 = i00 & n787;
  assign n793 = n760 & n792;
  assign n794 = ~n791 & ~n793;
  assign n795 = ~i04 & ~n794;
  assign n796 = ~n783 & ~n795;
  assign n797 = i03 & ~n796;
  assign n798 = ~i06 & n13;
  assign n799 = i06 & n14;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~i05 & ~n800;
  assign n802 = i05 & i06;
  assign n803 = n298 & n802;
  assign n804 = ~n801 & ~n803;
  assign n805 = i00 & ~n804;
  assign n806 = ~i06 & n298;
  assign n807 = n774 & n806;
  assign n808 = ~n805 & ~n807;
  assign n809 = i07 & ~n808;
  assign n810 = i04 & n809;
  assign n811 = ~i03 & n810;
  assign n812 = ~n797 & ~n811;
  assign n813 = i01 & ~n812;
  assign n814 = ~n767 & ~n813;
  assign n815 = ~n723 & ~n814;
  assign n816 = ~i02 & n98;
  assign n817 = i02 & n101;
  assign n818 = ~n816 & ~n817;
  assign n819 = i06 & ~n329;
  assign n820 = i00 & n819;
  assign n821 = ~i00 & i05;
  assign n822 = ~i06 & ~i09;
  assign n823 = n821 & n822;
  assign n824 = ~n820 & ~n823;
  assign n825 = ~i03 & ~n824;
  assign n826 = ~i06 & i09;
  assign n827 = ~i05 & n826;
  assign n828 = n75 & n827;
  assign n829 = ~n825 & ~n828;
  assign n830 = ~i10 & ~n829;
  assign n831 = i06 & ~i09;
  assign n832 = ~n826 & ~n831;
  assign n833 = i10 & ~n832;
  assign n834 = ~i05 & n833;
  assign n835 = ~i03 & n834;
  assign n836 = i00 & n835;
  assign n837 = ~n830 & ~n836;
  assign n838 = ~i01 & ~n837;
  assign n839 = i06 & n300;
  assign n840 = ~n806 & ~n839;
  assign n841 = ~i05 & ~n840;
  assign n842 = i03 & n841;
  assign n843 = i01 & n842;
  assign n844 = i00 & n843;
  assign n845 = ~n838 & ~n844;
  assign n846 = ~i07 & ~n845;
  assign n847 = n372 & n590;
  assign n848 = n366 & n473;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~i03 & ~n849;
  assign n851 = ~i00 & n850;
  assign n852 = i00 & n681;
  assign n853 = i05 & n465;
  assign n854 = n852 & n853;
  assign n855 = ~n851 & ~n854;
  assign n856 = ~i09 & ~n855;
  assign n857 = i07 & n856;
  assign n858 = ~n846 & ~n857;
  assign n859 = ~n818 & ~n858;
  assign n860 = i04 & i09;
  assign n861 = ~i04 & ~i09;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~i05 & i08;
  assign n864 = i05 & ~i08;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~i10 & ~n865;
  assign n867 = ~i07 & n866;
  assign n868 = i02 & n867;
  assign n869 = i05 & n342;
  assign n870 = ~i02 & n869;
  assign n871 = ~n868 & ~n870;
  assign n872 = i03 & ~n871;
  assign n873 = ~i03 & ~i05;
  assign n874 = i02 & n873;
  assign n875 = ~i07 & n493;
  assign n876 = n874 & n875;
  assign n877 = ~n872 & ~n876;
  assign n878 = ~i00 & ~n877;
  assign n879 = i07 & n479;
  assign n880 = ~i07 & n481;
  assign n881 = ~n879 & ~n880;
  assign n882 = i05 & ~n881;
  assign n883 = ~i03 & n882;
  assign n884 = n488 & n735;
  assign n885 = ~n883 & ~n884;
  assign n886 = i02 & ~n885;
  assign n887 = i00 & n886;
  assign n888 = ~n878 & ~n887;
  assign n889 = ~i06 & ~n888;
  assign n890 = i02 & n380;
  assign n891 = i05 & ~i07;
  assign n892 = ~i02 & n891;
  assign n893 = ~n890 & ~n892;
  assign n894 = i08 & ~n893;
  assign n895 = ~i03 & n894;
  assign n896 = i00 & n895;
  assign n897 = ~i00 & n564;
  assign n898 = i05 & n33;
  assign n899 = n897 & n898;
  assign n900 = ~n896 & ~n899;
  assign n901 = i10 & ~n900;
  assign n902 = i06 & n901;
  assign n903 = ~n889 & ~n902;
  assign n904 = ~i01 & ~n903;
  assign n905 = ~i05 & n232;
  assign n906 = ~n898 & ~n905;
  assign n907 = i10 & ~n906;
  assign n908 = i03 & n907;
  assign n909 = i00 & n908;
  assign n910 = ~n380 & ~n891;
  assign n911 = ~i10 & ~n910;
  assign n912 = i08 & n911;
  assign n913 = ~i03 & n912;
  assign n914 = ~i00 & n913;
  assign n915 = ~n909 & ~n914;
  assign n916 = i06 & ~n915;
  assign n917 = ~i00 & n735;
  assign n918 = n149 & n481;
  assign n919 = n917 & n918;
  assign n920 = ~n916 & ~n919;
  assign n921 = i02 & ~n920;
  assign n922 = n305 & n754;
  assign n923 = n148 & n487;
  assign n924 = n922 & n923;
  assign n925 = ~n921 & ~n924;
  assign n926 = i01 & ~n925;
  assign n927 = ~n904 & ~n926;
  assign n928 = ~n862 & ~n927;
  assign n929 = ~n784 & ~n787;
  assign n930 = i03 & ~n929;
  assign n931 = ~i03 & n787;
  assign n932 = ~n930 & ~n931;
  assign n933 = i09 & ~n932;
  assign n934 = ~i04 & n933;
  assign n935 = i05 & n831;
  assign n936 = n235 & n935;
  assign n937 = ~n934 & ~n936;
  assign n938 = ~i10 & ~n937;
  assign n939 = i04 & ~i05;
  assign n940 = i03 & n939;
  assign n941 = i06 & n13;
  assign n942 = n940 & n941;
  assign n943 = ~n938 & ~n942;
  assign n944 = ~i07 & ~n943;
  assign n945 = i05 & n298;
  assign n946 = ~i05 & n300;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~i04 & ~n947;
  assign n949 = n13 & n939;
  assign n950 = ~n948 & ~n949;
  assign n951 = i07 & ~n950;
  assign n952 = i06 & n951;
  assign n953 = i03 & n952;
  assign n954 = ~n944 & ~n953;
  assign n955 = i00 & ~n954;
  assign n956 = ~i04 & i05;
  assign n957 = n616 & n956;
  assign n958 = i07 & ~i10;
  assign n959 = n939 & n958;
  assign n960 = ~n957 & ~n959;
  assign n961 = i03 & ~n960;
  assign n962 = n235 & n869;
  assign n963 = ~n961 & ~n962;
  assign n964 = i09 & ~n963;
  assign n965 = i06 & n964;
  assign n966 = ~i00 & n965;
  assign n967 = ~n955 & ~n966;
  assign n968 = i01 & ~n967;
  assign n969 = n380 & n414;
  assign n970 = n606 & n891;
  assign n971 = ~n969 & ~n970;
  assign n972 = ~n357 & ~n971;
  assign n973 = ~i04 & ~i05;
  assign n974 = ~i00 & n973;
  assign n975 = n377 & n974;
  assign n976 = ~n972 & ~n975;
  assign n977 = i06 & ~n976;
  assign n978 = ~i00 & n939;
  assign n979 = n24 & n300;
  assign n980 = n978 & n979;
  assign n981 = ~n977 & ~n980;
  assign n982 = i03 & ~n981;
  assign n983 = ~i05 & n343;
  assign n984 = ~n869 & ~n983;
  assign n985 = ~i09 & ~n984;
  assign n986 = ~i06 & n985;
  assign n987 = i04 & n986;
  assign n988 = ~i03 & n987;
  assign n989 = ~i00 & n988;
  assign n990 = ~n982 & ~n989;
  assign n991 = ~i01 & ~n990;
  assign n992 = ~n968 & ~n991;
  assign n993 = i02 & ~n992;
  assign n994 = i03 & ~i06;
  assign n995 = ~n202 & ~n994;
  assign n996 = i09 & ~n995;
  assign n997 = ~i04 & n996;
  assign n998 = i00 & n997;
  assign n999 = i04 & n822;
  assign n1000 = n75 & n999;
  assign n1001 = ~n998 & ~n1000;
  assign n1002 = i05 & ~n1001;
  assign n1003 = i06 & i09;
  assign n1004 = i03 & n1003;
  assign n1005 = ~i03 & n822;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~i05 & ~n1006;
  assign n1008 = i04 & n1007;
  assign n1009 = ~i00 & n1008;
  assign n1010 = ~n1002 & ~n1009;
  assign n1011 = ~i01 & ~n1010;
  assign n1012 = n107 & n784;
  assign n1013 = n110 & n787;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = i09 & ~n1014;
  assign n1016 = i01 & n1015;
  assign n1017 = ~i00 & n1016;
  assign n1018 = ~n1011 & ~n1017;
  assign n1019 = ~i07 & ~n1018;
  assign n1020 = ~i01 & n1003;
  assign n1021 = i01 & n822;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~i03 & ~n1022;
  assign n1024 = ~i00 & n1023;
  assign n1025 = i00 & i01;
  assign n1026 = n1004 & n1025;
  assign n1027 = ~n1024 & ~n1026;
  assign n1028 = i07 & ~n1027;
  assign n1029 = ~i05 & n1028;
  assign n1030 = ~i04 & n1029;
  assign n1031 = ~n1019 & ~n1030;
  assign n1032 = i10 & ~n1031;
  assign n1033 = ~i06 & n737;
  assign n1034 = n42 & n1033;
  assign n1035 = i06 & n336;
  assign n1036 = n43 & n1035;
  assign n1037 = ~n1034 & ~n1036;
  assign n1038 = ~i00 & ~n1037;
  assign n1039 = i00 & n42;
  assign n1040 = i06 & n726;
  assign n1041 = n1039 & n1040;
  assign n1042 = ~n1038 & ~n1041;
  assign n1043 = ~i05 & ~n1042;
  assign n1044 = ~i04 & i09;
  assign n1045 = i04 & ~i09;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = i07 & ~n1046;
  assign n1048 = i06 & n1047;
  assign n1049 = i05 & n1048;
  assign n1050 = i01 & n1049;
  assign n1051 = i00 & n1050;
  assign n1052 = ~n1043 & ~n1051;
  assign n1053 = ~i10 & ~n1052;
  assign n1054 = i03 & n1053;
  assign n1055 = ~n1032 & ~n1054;
  assign n1056 = ~i02 & ~n1055;
  assign n1057 = ~n993 & ~n1056;
  assign n1058 = ~i08 & i09;
  assign n1059 = ~i07 & n1058;
  assign n1060 = n645 & n1059;
  assign n1061 = i08 & ~i09;
  assign n1062 = i07 & n1061;
  assign n1063 = n203 & n1062;
  assign n1064 = ~n1060 & ~n1063;
  assign n1065 = i01 & i10;
  assign n1066 = ~i01 & ~i10;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = i05 & ~n1067;
  assign n1069 = i03 & n1068;
  assign n1070 = i02 & n1069;
  assign n1071 = i00 & n1070;
  assign n1072 = ~i00 & n464;
  assign n1073 = ~i03 & n769;
  assign n1074 = n1072 & n1073;
  assign n1075 = ~n1071 & ~n1074;
  assign n1076 = ~n1064 & ~n1075;
  assign n1077 = ~i04 & n730;
  assign n1078 = i04 & n726;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = i02 & ~i03;
  assign n1081 = ~i01 & n1080;
  assign n1082 = ~i05 & n108;
  assign n1083 = n1081 & n1082;
  assign n1084 = i01 & n510;
  assign n1085 = i05 & n111;
  assign n1086 = n1084 & n1085;
  assign n1087 = ~n1083 & ~n1086;
  assign n1088 = i00 & ~n1087;
  assign n1089 = i03 & i05;
  assign n1090 = n111 & n1089;
  assign n1091 = n1072 & n1090;
  assign n1092 = ~n1088 & ~n1091;
  assign n1093 = i10 & ~n1092;
  assign n1094 = ~i00 & ~i01;
  assign n1095 = n510 & n1094;
  assign n1096 = n493 & n787;
  assign n1097 = n1095 & n1096;
  assign n1098 = ~n1093 & ~n1097;
  assign n1099 = ~n1079 & ~n1098;
  assign n1100 = i02 & n232;
  assign n1101 = ~i02 & n33;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = ~i03 & n298;
  assign n1104 = i03 & n300;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~i05 & ~n1105;
  assign n1107 = i00 & n1106;
  assign n1108 = i05 & n13;
  assign n1109 = n75 & n1108;
  assign n1110 = ~n1107 & ~n1109;
  assign n1111 = i06 & ~n1110;
  assign n1112 = i04 & n1111;
  assign n1113 = ~i06 & ~n357;
  assign n1114 = i05 & n1113;
  assign n1115 = ~i04 & n1114;
  assign n1116 = i03 & n1115;
  assign n1117 = ~i00 & n1116;
  assign n1118 = ~n1112 & ~n1117;
  assign n1119 = i01 & ~n1118;
  assign n1120 = ~n460 & ~n465;
  assign n1121 = i05 & ~n1120;
  assign n1122 = ~i05 & n473;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~i09 & ~n1123;
  assign n1125 = i00 & n1124;
  assign n1126 = n774 & n799;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = i04 & ~n1127;
  assign n1129 = ~i03 & n1128;
  assign n1130 = ~i01 & n1129;
  assign n1131 = ~n1119 & ~n1130;
  assign n1132 = ~n1102 & ~n1131;
  assign n1133 = n100 & n826;
  assign n1134 = n97 & n831;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = i00 & ~n1135;
  assign n1137 = i03 & n831;
  assign n1138 = n362 & n1137;
  assign n1139 = ~n1136 & ~n1138;
  assign n1140 = ~i08 & ~n1139;
  assign n1141 = i01 & n826;
  assign n1142 = ~i01 & n831;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = i08 & ~n1143;
  assign n1145 = ~i03 & n1144;
  assign n1146 = ~i00 & n1145;
  assign n1147 = ~n1140 & ~n1146;
  assign n1148 = ~i10 & ~n1147;
  assign n1149 = n108 & n298;
  assign n1150 = n682 & n1149;
  assign n1151 = ~n1148 & ~n1150;
  assign n1152 = i05 & ~n1151;
  assign n1153 = n362 & n873;
  assign n1154 = n111 & n298;
  assign n1155 = n1153 & n1154;
  assign n1156 = ~n1152 & ~n1155;
  assign n1157 = n487 & n821;
  assign n1158 = i00 & ~i05;
  assign n1159 = n493 & n1158;
  assign n1160 = ~n1157 & ~n1159;
  assign n1161 = i02 & ~n1160;
  assign n1162 = ~n479 & ~n481;
  assign n1163 = i00 & ~n1162;
  assign n1164 = ~i00 & n493;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~i05 & ~n1165;
  assign n1167 = n481 & n821;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~i02 & ~n1168;
  assign n1170 = ~n1161 & ~n1169;
  assign n1171 = i01 & ~n1170;
  assign n1172 = ~i05 & i10;
  assign n1173 = i05 & ~i10;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = i00 & ~n1174;
  assign n1176 = ~i00 & n1173;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = ~i02 & ~n1177;
  assign n1179 = n433 & n769;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = ~i08 & ~n1180;
  assign n1182 = i08 & ~n1174;
  assign n1183 = i02 & n1182;
  assign n1184 = i00 & n1183;
  assign n1185 = ~n1181 & ~n1184;
  assign n1186 = ~i01 & ~n1185;
  assign n1187 = ~n1171 & ~n1186;
  assign n1188 = ~i09 & ~n1187;
  assign n1189 = ~i00 & ~i10;
  assign n1190 = i00 & n636;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~i02 & ~n1191;
  assign n1193 = i00 & n471;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = i08 & ~n1194;
  assign n1196 = i00 & ~i01;
  assign n1197 = i02 & n481;
  assign n1198 = n1196 & n1197;
  assign n1199 = ~n1195 & ~n1198;
  assign n1200 = ~i05 & ~n1199;
  assign n1201 = i00 & n310;
  assign n1202 = i05 & n479;
  assign n1203 = n1201 & n1202;
  assign n1204 = ~n1200 & ~n1203;
  assign n1205 = i09 & ~n1204;
  assign n1206 = ~n1188 & ~n1205;
  assign n1207 = ~i06 & ~n1206;
  assign n1208 = i02 & i09;
  assign n1209 = ~i02 & ~i09;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~i01 & ~n1162;
  assign n1212 = i00 & n1211;
  assign n1213 = n362 & n487;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1210 & ~n1214;
  assign n1216 = ~i01 & i08;
  assign n1217 = ~i00 & n1216;
  assign n1218 = i01 & ~i08;
  assign n1219 = i00 & n1218;
  assign n1220 = ~n1217 & ~n1219;
  assign n1221 = i10 & ~n1220;
  assign n1222 = ~i09 & n1221;
  assign n1223 = ~i02 & n1222;
  assign n1224 = ~n1215 & ~n1223;
  assign n1225 = ~i05 & ~n1224;
  assign n1226 = ~i02 & ~n1162;
  assign n1227 = i01 & n1226;
  assign n1228 = n310 & n479;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~i00 & ~n1229;
  assign n1231 = ~i02 & n487;
  assign n1232 = n1196 & n1231;
  assign n1233 = ~n1230 & ~n1232;
  assign n1234 = i09 & ~n1233;
  assign n1235 = i05 & n1234;
  assign n1236 = ~n1225 & ~n1235;
  assign n1237 = i06 & ~n1236;
  assign n1238 = ~n1207 & ~n1237;
  assign n1239 = i03 & ~n1238;
  assign n1240 = n45 & n298;
  assign n1241 = n48 & n300;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~i02 & ~n1242;
  assign n1244 = i08 & n298;
  assign n1245 = ~i08 & n300;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~i06 & ~n1246;
  assign n1248 = ~n1154 & ~n1247;
  assign n1249 = i02 & ~n1248;
  assign n1250 = ~n1243 & ~n1249;
  assign n1251 = i00 & ~n1250;
  assign n1252 = i09 & ~n298;
  assign n1253 = ~i08 & ~n1252;
  assign n1254 = ~i06 & n1253;
  assign n1255 = n13 & n48;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = i02 & ~n1256;
  assign n1258 = ~i00 & n1257;
  assign n1259 = ~n1251 & ~n1258;
  assign n1260 = ~i01 & ~n1259;
  assign n1261 = i00 & i10;
  assign n1262 = ~i00 & n473;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = i08 & ~n1263;
  assign n1265 = n487 & n725;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = i09 & ~n1266;
  assign n1268 = i00 & i06;
  assign n1269 = ~i08 & n13;
  assign n1270 = n1268 & n1269;
  assign n1271 = ~n1267 & ~n1270;
  assign n1272 = ~i02 & ~n1271;
  assign n1273 = i01 & n1272;
  assign n1274 = ~n1260 & ~n1273;
  assign n1275 = ~i05 & ~n1274;
  assign n1276 = i00 & ~n691;
  assign n1277 = ~n1094 & ~n1276;
  assign n1278 = i09 & ~n1277;
  assign n1279 = ~i00 & n822;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~i10 & ~n1280;
  assign n1282 = n806 & n1094;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~i08 & ~n1283;
  assign n1285 = ~i01 & i06;
  assign n1286 = i00 & n1285;
  assign n1287 = n1244 & n1286;
  assign n1288 = ~n1284 & ~n1287;
  assign n1289 = ~i02 & ~n1288;
  assign n1290 = n45 & n300;
  assign n1291 = n1193 & n1290;
  assign n1292 = ~n1289 & ~n1291;
  assign n1293 = i05 & ~n1292;
  assign n1294 = ~n1275 & ~n1293;
  assign n1295 = ~i03 & ~n1294;
  assign n1296 = ~n1239 & ~n1295;
  assign n1297 = n1156 & n1296;
  assign n1298 = i07 & ~n1297;
  assign n1299 = ~i05 & n481;
  assign n1300 = ~n1202 & ~n1299;
  assign n1301 = ~i03 & ~n1300;
  assign n1302 = i02 & n1301;
  assign n1303 = i05 & n481;
  assign n1304 = ~n863 & ~n1303;
  assign n1305 = i03 & ~n1304;
  assign n1306 = ~i02 & n1305;
  assign n1307 = ~n1302 & ~n1306;
  assign n1308 = i01 & ~n1307;
  assign n1309 = i02 & ~n770;
  assign n1310 = ~i02 & ~n1174;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = i08 & ~n1311;
  assign n1313 = i03 & n1312;
  assign n1314 = i05 & n487;
  assign n1315 = n1080 & n1314;
  assign n1316 = ~n1313 & ~n1315;
  assign n1317 = ~i01 & ~n1316;
  assign n1318 = ~n1308 & ~n1317;
  assign n1319 = i09 & ~n1318;
  assign n1320 = i02 & i05;
  assign n1321 = ~i02 & ~i05;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = i01 & ~i03;
  assign n1324 = ~n681 & ~n1323;
  assign n1325 = ~n1322 & ~n1324;
  assign n1326 = ~i08 & n1325;
  assign n1327 = i05 & i08;
  assign n1328 = ~i03 & n1327;
  assign n1329 = ~i01 & n1328;
  assign n1330 = ~n1326 & ~n1329;
  assign n1331 = ~i10 & ~n1330;
  assign n1332 = ~i01 & n551;
  assign n1333 = n1314 & n1332;
  assign n1334 = ~n1331 & ~n1333;
  assign n1335 = ~i09 & ~n1334;
  assign n1336 = ~n1319 & ~n1335;
  assign n1337 = i06 & ~n1336;
  assign n1338 = i09 & ~n1174;
  assign n1339 = ~i01 & n1338;
  assign n1340 = n300 & n372;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = i02 & ~n1341;
  assign n1343 = ~i10 & ~n329;
  assign n1344 = ~i02 & n1343;
  assign n1345 = i01 & n1344;
  assign n1346 = ~n1342 & ~n1345;
  assign n1347 = ~i03 & ~n1346;
  assign n1348 = ~i01 & n327;
  assign n1349 = ~n386 & ~n1348;
  assign n1350 = i10 & ~n1349;
  assign n1351 = ~i02 & n1350;
  assign n1352 = n471 & n946;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = i03 & ~n1353;
  assign n1355 = ~n1347 & ~n1354;
  assign n1356 = i08 & ~n1355;
  assign n1357 = i03 & i10;
  assign n1358 = ~i03 & n300;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~i05 & ~n1359;
  assign n1361 = ~i01 & n1360;
  assign n1362 = n312 & n1323;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = ~i08 & ~n1363;
  assign n1365 = ~i02 & n1364;
  assign n1366 = ~n1356 & ~n1365;
  assign n1367 = ~i06 & ~n1366;
  assign n1368 = ~n1337 & ~n1367;
  assign n1369 = ~i00 & ~n1368;
  assign n1370 = n108 & n1320;
  assign n1371 = n111 & n1321;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = i03 & i09;
  assign n1374 = ~i03 & ~i09;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = ~n1372 & ~n1375;
  assign n1377 = i02 & ~i09;
  assign n1378 = i02 & ~n1377;
  assign n1379 = i08 & ~n1378;
  assign n1380 = ~i06 & n1379;
  assign n1381 = i05 & n1380;
  assign n1382 = i03 & n1381;
  assign n1383 = ~n1376 & ~n1382;
  assign n1384 = ~i01 & ~n1383;
  assign n1385 = ~i02 & i05;
  assign n1386 = i06 & n1058;
  assign n1387 = n1385 & n1386;
  assign n1388 = i02 & ~i05;
  assign n1389 = ~i06 & n1061;
  assign n1390 = n1388 & n1389;
  assign n1391 = ~n1387 & ~n1390;
  assign n1392 = i03 & ~n1391;
  assign n1393 = ~i09 & ~n865;
  assign n1394 = i02 & n1393;
  assign n1395 = n1058 & n1385;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~i06 & ~n1396;
  assign n1398 = ~i05 & n1058;
  assign n1399 = i05 & n1061;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = i06 & ~n1400;
  assign n1402 = ~i02 & n1401;
  assign n1403 = ~n1397 & ~n1402;
  assign n1404 = ~i03 & ~n1403;
  assign n1405 = ~n1392 & ~n1404;
  assign n1406 = i01 & ~n1405;
  assign n1407 = ~n1384 & ~n1406;
  assign n1408 = ~i10 & ~n1407;
  assign n1409 = i02 & n202;
  assign n1410 = ~i02 & n994;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~i05 & ~n1411;
  assign n1413 = i01 & n1412;
  assign n1414 = ~i02 & ~i06;
  assign n1415 = ~i02 & ~n1414;
  assign n1416 = i05 & ~n1415;
  assign n1417 = ~i03 & n1416;
  assign n1418 = ~i01 & n1417;
  assign n1419 = ~n1413 & ~n1418;
  assign n1420 = ~i09 & ~n1419;
  assign n1421 = i01 & ~n457;
  assign n1422 = ~i01 & n403;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = i09 & ~n1423;
  assign n1425 = ~i05 & n1424;
  assign n1426 = i03 & n1425;
  assign n1427 = ~n1420 & ~n1426;
  assign n1428 = i08 & ~n1427;
  assign n1429 = ~i01 & n510;
  assign n1430 = ~i08 & ~i09;
  assign n1431 = n802 & n1430;
  assign n1432 = n1429 & n1431;
  assign n1433 = ~n1428 & ~n1432;
  assign n1434 = i10 & ~n1433;
  assign n1435 = ~n1408 & ~n1434;
  assign n1436 = i00 & ~n1435;
  assign n1437 = ~n1369 & ~n1436;
  assign n1438 = ~i07 & ~n1437;
  assign n1439 = ~n1298 & ~n1438;
  assign n1440 = ~i04 & ~n1439;
  assign n1441 = i01 & i09;
  assign n1442 = ~i01 & ~i09;
  assign n1443 = ~n1441 & ~n1442;
  assign n1444 = ~i02 & ~n1443;
  assign n1445 = i00 & n1444;
  assign n1446 = ~i01 & i09;
  assign n1447 = i01 & ~i09;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = i02 & ~n1448;
  assign n1450 = ~i00 & n1449;
  assign n1451 = ~n1445 & ~n1450;
  assign n1452 = i05 & ~n1451;
  assign n1453 = ~i05 & i09;
  assign n1454 = ~i01 & n1453;
  assign n1455 = i00 & n1454;
  assign n1456 = ~n1452 & ~n1455;
  assign n1457 = ~i03 & ~n1456;
  assign n1458 = ~n310 & ~n464;
  assign n1459 = ~i00 & ~n1458;
  assign n1460 = ~n1201 & ~n1459;
  assign n1461 = i09 & ~n1460;
  assign n1462 = ~i05 & n1461;
  assign n1463 = i03 & n1462;
  assign n1464 = ~n1457 & ~n1463;
  assign n1465 = i07 & ~n1464;
  assign n1466 = i05 & ~i09;
  assign n1467 = ~n1453 & ~n1466;
  assign n1468 = i00 & n510;
  assign n1469 = ~i00 & n1080;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = ~n1467 & ~n1470;
  assign n1472 = ~i09 & ~n76;
  assign n1473 = i05 & n1472;
  assign n1474 = i02 & n1473;
  assign n1475 = ~n1471 & ~n1474;
  assign n1476 = ~i01 & ~n1475;
  assign n1477 = ~i02 & ~n510;
  assign n1478 = ~i05 & ~n1477;
  assign n1479 = ~i02 & n754;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = ~i09 & ~n1480;
  assign n1482 = i01 & n1481;
  assign n1483 = ~i00 & n1482;
  assign n1484 = ~n1476 & ~n1483;
  assign n1485 = ~i07 & ~n1484;
  assign n1486 = ~n1465 & ~n1485;
  assign n1487 = ~i08 & ~n1486;
  assign n1488 = n327 & n551;
  assign n1489 = n328 & n564;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~i01 & ~n1490;
  assign n1492 = i05 & ~n1375;
  assign n1493 = ~i02 & n1492;
  assign n1494 = n1080 & n1453;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = i01 & ~n1495;
  assign n1497 = ~n1491 & ~n1496;
  assign n1498 = i07 & ~n1497;
  assign n1499 = ~i01 & n873;
  assign n1500 = n100 & n1466;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = ~i07 & ~n1501;
  assign n1503 = i02 & n1502;
  assign n1504 = ~n1498 & ~n1503;
  assign n1505 = i00 & ~n1504;
  assign n1506 = ~i03 & n380;
  assign n1507 = i03 & n891;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = i01 & ~n1508;
  assign n1510 = n97 & n354;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~i09 & ~n1511;
  assign n1513 = ~i05 & n730;
  assign n1514 = n681 & n1513;
  assign n1515 = ~n1512 & ~n1514;
  assign n1516 = i02 & ~n1515;
  assign n1517 = ~i05 & n737;
  assign n1518 = n1332 & n1517;
  assign n1519 = ~n1516 & ~n1518;
  assign n1520 = ~i00 & ~n1519;
  assign n1521 = ~n1505 & ~n1520;
  assign n1522 = i08 & ~n1521;
  assign n1523 = ~n1487 & ~n1522;
  assign n1524 = i06 & ~n1523;
  assign n1525 = i03 & n415;
  assign n1526 = ~i03 & n1430;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = i00 & ~n1527;
  assign n1529 = ~i03 & i09;
  assign n1530 = i03 & ~i09;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = i08 & ~n1531;
  assign n1533 = ~i00 & n1532;
  assign n1534 = ~n1528 & ~n1533;
  assign n1535 = ~i02 & ~n1534;
  assign n1536 = ~n1058 & ~n1061;
  assign n1537 = i03 & ~n1536;
  assign n1538 = i02 & n1537;
  assign n1539 = ~i00 & n1538;
  assign n1540 = ~n1535 & ~n1539;
  assign n1541 = i07 & ~n1540;
  assign n1542 = ~i08 & ~n1210;
  assign n1543 = i00 & n1542;
  assign n1544 = n433 & n1061;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~i03 & ~n1545;
  assign n1547 = i03 & n1061;
  assign n1548 = n433 & n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign n1550 = ~i07 & ~n1549;
  assign n1551 = ~n1541 & ~n1550;
  assign n1552 = i01 & ~n1551;
  assign n1553 = ~n510 & ~n1080;
  assign n1554 = i00 & ~n1553;
  assign n1555 = ~n1469 & ~n1554;
  assign n1556 = ~i08 & ~n1555;
  assign n1557 = i07 & n1556;
  assign n1558 = i03 & n17;
  assign n1559 = n305 & n1558;
  assign n1560 = ~n1557 & ~n1559;
  assign n1561 = ~i09 & ~n1560;
  assign n1562 = i07 & n1058;
  assign n1563 = ~i02 & n1562;
  assign n1564 = i00 & n1563;
  assign n1565 = ~n1561 & ~n1564;
  assign n1566 = ~i01 & ~n1565;
  assign n1567 = ~n1552 & ~n1566;
  assign n1568 = ~i05 & ~n1567;
  assign n1569 = ~n415 & ~n1430;
  assign n1570 = n119 & n1196;
  assign n1571 = n127 & n362;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = ~n1569 & ~n1572;
  assign n1574 = i03 & n726;
  assign n1575 = ~n1529 & ~n1574;
  assign n1576 = ~i08 & ~n1575;
  assign n1577 = i01 & n1576;
  assign n1578 = i00 & n1577;
  assign n1579 = ~i00 & n97;
  assign n1580 = n1062 & n1579;
  assign n1581 = ~n1578 & ~n1580;
  assign n1582 = ~n1573 & n1581;
  assign n1583 = ~i02 & ~n1582;
  assign n1584 = n116 & n1430;
  assign n1585 = n1193 & n1584;
  assign n1586 = ~n1583 & ~n1585;
  assign n1587 = i05 & ~n1586;
  assign n1588 = ~n1568 & ~n1587;
  assign n1589 = ~i06 & ~n1588;
  assign n1590 = ~n1524 & ~n1589;
  assign n1591 = ~i10 & ~n1590;
  assign n1592 = n310 & n1089;
  assign n1593 = n464 & n873;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~i07 & ~n1594;
  assign n1596 = i00 & n1595;
  assign n1597 = n472 & n1506;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = i08 & ~n1598;
  assign n1600 = ~i01 & ~i02;
  assign n1601 = i00 & n1600;
  assign n1602 = n20 & n1089;
  assign n1603 = n1601 & n1602;
  assign n1604 = ~n1599 & ~n1603;
  assign n1605 = i07 & n415;
  assign n1606 = n100 & n1605;
  assign n1607 = ~i07 & n1430;
  assign n1608 = n97 & n1607;
  assign n1609 = ~n1606 & ~n1608;
  assign n1610 = i00 & ~n1609;
  assign n1611 = ~n33 & ~n232;
  assign n1612 = i01 & ~n1611;
  assign n1613 = ~i01 & ~n456;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = i09 & ~n1614;
  assign n1616 = n699 & n1061;
  assign n1617 = ~n1615 & ~n1616;
  assign n1618 = i03 & ~n1617;
  assign n1619 = n1059 & n1323;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~i00 & ~n1620;
  assign n1622 = ~n1610 & ~n1621;
  assign n1623 = ~i05 & ~n1622;
  assign n1624 = ~i09 & ~n548;
  assign n1625 = ~i07 & n1624;
  assign n1626 = i05 & n1625;
  assign n1627 = ~i01 & n1626;
  assign n1628 = ~i00 & n1627;
  assign n1629 = ~n1623 & ~n1628;
  assign n1630 = i02 & ~n1629;
  assign n1631 = n737 & n873;
  assign n1632 = n336 & n1089;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = i00 & ~n1633;
  assign n1635 = i05 & n737;
  assign n1636 = n123 & n1635;
  assign n1637 = ~n1634 & ~n1636;
  assign n1638 = i08 & ~n1637;
  assign n1639 = ~n873 & ~n1089;
  assign n1640 = ~i09 & ~n1639;
  assign n1641 = ~i08 & n1640;
  assign n1642 = i07 & n1641;
  assign n1643 = ~i00 & n1642;
  assign n1644 = ~n1638 & ~n1643;
  assign n1645 = ~i02 & ~n1644;
  assign n1646 = ~i01 & n1645;
  assign n1647 = ~n1630 & ~n1646;
  assign n1648 = n1604 & n1647;
  assign n1649 = ~i06 & ~n1648;
  assign n1650 = ~i07 & n1061;
  assign n1651 = ~n1562 & ~n1650;
  assign n1652 = i02 & ~n1651;
  assign n1653 = ~i02 & n1058;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~i05 & ~n1654;
  assign n1656 = n1062 & n1320;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = ~i00 & ~n1657;
  assign n1659 = n200 & n1058;
  assign n1660 = ~n1652 & ~n1659;
  assign n1661 = i05 & ~n1660;
  assign n1662 = n1321 & n1562;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = i00 & ~n1663;
  assign n1665 = ~n1658 & ~n1664;
  assign n1666 = ~i01 & ~n1665;
  assign n1667 = i02 & n730;
  assign n1668 = ~i02 & n726;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = i00 & ~n1669;
  assign n1671 = ~n726 & ~n730;
  assign n1672 = i02 & ~n1671;
  assign n1673 = ~i00 & n1672;
  assign n1674 = ~n1670 & ~n1673;
  assign n1675 = ~i08 & ~n1674;
  assign n1676 = ~i05 & n1675;
  assign n1677 = i01 & n1676;
  assign n1678 = ~n1666 & ~n1677;
  assign n1679 = ~i03 & ~n1678;
  assign n1680 = i00 & i02;
  assign n1681 = n415 & n1680;
  assign n1682 = n305 & n1430;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n356 & ~n1683;
  assign n1685 = n199 & n1061;
  assign n1686 = ~n1659 & ~n1685;
  assign n1687 = ~i05 & ~n1686;
  assign n1688 = i00 & n1687;
  assign n1689 = ~n176 & ~n320;
  assign n1690 = i09 & ~n1689;
  assign n1691 = i08 & n1690;
  assign n1692 = i05 & n1691;
  assign n1693 = ~i00 & n1692;
  assign n1694 = ~n1688 & ~n1693;
  assign n1695 = ~n1684 & n1694;
  assign n1696 = i03 & ~n1695;
  assign n1697 = ~i01 & n1696;
  assign n1698 = ~n1679 & ~n1697;
  assign n1699 = i06 & ~n1698;
  assign n1700 = ~n1649 & ~n1699;
  assign n1701 = i10 & ~n1700;
  assign n1702 = ~n1591 & ~n1701;
  assign n1703 = i04 & ~n1702;
  assign n1704 = ~n1440 & ~n1703;
  assign n1705 = ~n1132 & n1704;
  assign n1706 = ~n1099 & n1705;
  assign n1707 = ~n1076 & n1706;
  assign n1708 = n1057 & n1707;
  assign n1709 = ~n928 & n1708;
  assign n1710 = ~n859 & n1709;
  assign n1711 = ~n815 & n1710;
  assign n1712 = n720 & n1711;
  assign n1713 = ~n395 & n1712;
  assign f = n295 | ~n1713;
endmodule


